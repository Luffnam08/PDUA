--------------------------------------------------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
--------------------------------------------------------------------------------------------------------------------------
ENTITY upROM IS
	GENERIC(A_Bits : INTEGER := 8;
			  W_Bits : INTEGER := 29);
   PORT(   clk    : IN  STD_LOGIC;
			  addr   : IN  STD_LOGIC_VECTOR(A_Bits-1 DOWNTO 0);
		     r_data : OUT STD_LOGIC_VECTOR(W_Bits-1 DOWNTO 0));
END ENTITY upROM;	
--------------------------------------------------------------------------------------------------------------------------
ARCHITECTURE RTL OF upROM IS
TYPE mem_type IS ARRAY (0 TO 2**A_Bits-1) OF STD_LOGIC_VECTOR(W_Bits-1 DOWNTO 0);
SIGNAL rom : mem_type := (
--FETCH-------------------------------------------------------------------------------------------------------------------
0   => b"00000000000000001000010000000", 1   => b"00000000000001011000010000000", 2   => b"00000000000000011000010000000",
3   => b"00000000000000011001010000000", 4   => b"01100000000000001000011000000", 5   => b"00000000000010001000010000000",
--MOV ACC, A--------------------------------------------------------------------------------------------------------------
8   => b"00000001111100001000011000000", 9   => b"10000001111110001000110000000",
--MOV A, ACC--------------------------------------------------------------------------------------------------------------
16  => b"00000011101100001000011000000", 17  => b"10000011101110001000110000000",
--MOV ACC, CTE------------------------------------------------------------------------------------------------------------
24  => b"00000000011100001000010000000", 25  => b"00000000011101011000010000000", 26  => b"00000000011100011000010000000",
27  => b"00000000011110011000010000000", 28  => b"01100000000000001000011000000", 29  => b"00000000000010001000110000000",
--MOV ACC, [DPTR]---------------------------------------------------------------------------------------------------------
32  => b"00000001011100001000010000000", 33  => b"00000001011101011000010000000", 34  => b"00000001011100011000011000000",
35  => b"00000001011110011000110000000",
--MOV DPTR, ACC-----------------------------------------------------------------------------------------------------------
40  => b"00000011101000001000011000000", 41  => b"10000011101010001000110000000",
--MOV [DPTR], ACC---------------------------------------------------------------------------------------------------------
48  => b"00000001000000001000010000000", 49  => b"00000001000001011000010000000", 50  => b"00000011100000101000011000000",
51  => b"10000011100000101010110000000",
--INV ACC-----------------------------------------------------------------------------------------------------------------
56  => b"00010011111100001000011000000", 57  => b"10010011111110001000110000000",
--AND ACC, A--------------------------------------------------------------------------------------------------------------
64  => b"00000000000000001000011000000", 65  => b"00000000000000001000110000000",
--ADD ACC, A--------------------------------------------------------------------------------------------------------------
72  => b"00100001111100001000011000000", 73  => b"10100001111110001000110000000",
--JMP CTE-----------------------------------------------------------------------------------------------------------------
80  => b"00000000000000000000000000000", 81  => b"00000000000000000000000000000", 82  => b"00000000000000000000000000000",
83  => b"00000000000000000000000000000", 84  => b"00000000000000000000000000000", 85  => b"00000000000000000000000000000",
86  => b"00000000000000000000000000000", 87  => b"00000000000000000000000000000",
--JZ CTE------------------------------------------------------------------------------------------------------------------
88  => b"00000000000000000000000000000", 89  => b"00000000000000000000000000000", 90  => b"00000000000000000000000000000",
91  => b"00000000000000000000000000000", 92  => b"00000000000000000000000000000", 93  => b"00000000000000000000000000000",
94  => b"00000000000000000000000000000", 95  => b"00000000000000000000000000000",
--JN CTE------------------------------------------------------------------------------------------------------------------
96  => b"00000000000000000000000000000", 97  => b"00000000000000000000000000000", 98  => b"00000000000000000000000000000",
99  => b"00000000000000000000000000000", 100 => b"00000000000000000000000000000", 101 => b"00000000000000000000000000000",
102 => b"00000000000000000000000000000", 103 => b"00000000000000000000000000000",
--JC CTE------------------------------------------------------------------------------------------------------------------
104 => b"00000000000000000000000000000", 105 => b"00000000000000000000000000000", 106 => b"00000000000000000000000000000",
107 => b"00000000000000000000000000000", 108 => b"00000000000000000000000000000", 109 => b"00000000000000000000000000000",
110 => b"00000000000000000000000000000", 111 => b"00000000000000000000000000000",
--CALL DIR----------------------------------------------------------------------------------------------------------------
112 => b"00000000000000000000000000000", 113 => b"00000000000000000000000000000", 114 => b"00000000000000000000000000000",
115 => b"00000000000000000000000000000", 116 => b"00000000000000000000000000000", 117 => b"00000000000000000000000000000",
118 => b"00000000000000000000000000000", 119 => b"00000000000000000000000000000",
--RET---------------------------------------------------------------------------------------------------------------------
120 => b"00000000000000000000000000000", 121 => b"00000000000000000000000000000", 122 => b"00000000000000000000000000000",
123 => b"00000000000000000000000000000", 124 => b"00000000000000000000000000000", 125 => b"00000000000000000000000000000",
126 => b"00000000000000000000000000000", 127 => b"00000000000000000000000000000",
--MOV DPTR, CTE-----------------------------------------------------------------------------------------------------------
128 => b"00000000001000001000010000000", 129 => b"00000000001001011000010000000", 130 => b"00000000001000011000010000000",
131 => b"00000000001010011000010000000", 132 => b"01100000000000001000011000000", 133 => b"00000000000010001000110000000",
--MOV A, [DPTR]-----------------------------------------------------------------------------------------------------------
136 => b"00000001001100001000010000000", 137 => b"00000001001101011000010000000", 138 => b"00000001001100011000011000000",
139 => b"00000001001110011000110000000",
--NEG ACC-----------------------------------------------------------------------------------------------------------------
144 => b"01110011111100001000011000000", 145 => b"11110011111110001000110000000",
--INC ACC-----------------------------------------------------------------------------------------------------------------
152 => b"01100011111100001000011000000", 153 => b"11100011111110001000110000000",
--DEC ACC-----------------------------------------------------------------------------------------------------------------
160 => b"01010011011100001000011000000", 161 => b"11010011011110001000110000000",
--OR ACC, A---------------------------------------------------------------------------------------------------------------
168 => b"00110001111100001000011000000", 169 => b"10110001111110001000110000000",
--XOR ACC, A--------------------------------------------------------------------------------------------------------------
176 => b"01000001111100001000011000000", 177 => b"11000001111110001000110000000",
--SLL ACC-----------------------------------------------------------------------------------------------------------------
184 => b"00001011111100001000011000000", 185 => b"10001011111110001000110000000",
--SLR ACC-----------------------------------------------------------------------------------------------------------------
192 => b"00000111111100001000011000000", 193 => b"10000111111110001000110000000",
--LSB ACC-----------------------------------------------------------------------------------------------------------------
200 => b"01110011010100001000010000000", 201 => b"01110011010110001000010000000", 202 => b"00100010111100001000011000000",
203 => b"10100010111110001000110000000",
--NAND ACC, A-------------------------------------------------------------------------------------------------------------
208 => b"00100001110100001000010000000", 209 => b"10100001110110001000010000000", 210 => b"00010010111100001000011000000",
211 => b"10010010111110001000110000000",
--HALT--------------------------------------------------------------------------------------------------------------------
216 => b"00000000000000001000111000000",
--------------------------------------------------------------------------------------------------------------------------
OTHERS => b"00000000000000000000000000000");
--------------------------------------------------------------------------------------------------------------------------
BEGIN
	write_process: PROCESS(clk)
	BEGIN	
		IF (RISING_EDGE(clk)) THEN
			r_data <= rom(TO_INTEGER(UNSIGNED(addr)));
		END IF;
	END PROCESS;
--------------------------------------------------------------------------------------------------------------------------
END ARCHITECTURE RTL;
--------------------------------------------------------------------------------------------------------------------------